class transaction;
  
  bit [7:0]instrMem [0:1023]; //Modified from 63 to 1023
  
endclass